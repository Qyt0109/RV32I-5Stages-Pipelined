module execute ();

endmodule
