module decode ();

endmodule
