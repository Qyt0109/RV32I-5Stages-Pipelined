module fetch (
    
);

endmodule
