module forward (
    
);
    
endmodule